module mux_3x1_16bit_tb ();
    reg [1:0] S;
    reg [15:0] A, B, C;
    wire [15:0] X;
    
    integer errors = 0;

    task Check;
        input [31:0] expect;
        if (expect[31:16] != expect[15:0]) begin
            $display("Got %d, expected %d", expect[31:16], expect[15:0]);
            errors = errors + 1;
        end
    endtask

    mux_3x1_16bit UUT (.A(A), .B(B), .C(C), .X(X), .S(S));

    initial begin
       #10
       S <= 2'b00; 
       A <= 16'd1; B <= 16'd2; C <= 16'd3;
       
       #10

       $display("Test saida A");
       S <= 2'b00;
       #10
       Check({X, A});
       #10

       $display("Test saida B");
       S = 2'b01;
       #10
       Check({X, B});
       #10

       $display("Test saida C");
       S = 2'b10;
       #10
       Check({X, C});
       #10

       $display("Errors: %d", errors);
       $finish;
       
    end
endmodule